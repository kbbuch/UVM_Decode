package decode_in_pkg;
  
    import uvm_pkg::*;
    
    /*****************TX VIEW***************/
    import questa_uvm_pkg::*;
    /*****************TX VIEW***************/
    
    `include "uvm_macros.svh"
  
    `include "src/decode_seq_item.svh"
    
    `include "src/decode_config.svh"
    `include "src/decode_coverage.svh"
    
    `include "src/decode_sequence.svh"
    `include "src/decode_sequencer.svh"
    `include "src/decode_driver.svh"
    `include "src/decode_monitor.svh"
    `include "src/decode_agent.svh"

endpackage
