package decode_test_pkg;
  
    import uvm_pkg::*;
   import decode_in_pkg::*; 
   import decode_out_pkg::*; 
   import uvmf_base_pkg_hdl::*;
	import uvmf_base_pkg::*;
    `include "uvm_macros.svh"
  
    `include "src/test_top.svh"

endpackage
